library verilog;
use verilog.vl_types.all;
entity uart_TB is
end uart_TB;
